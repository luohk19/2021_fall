library verilog;
use verilog.vl_types.all;
entity scanning_tb is
end scanning_tb;
