library verilog;
use verilog.vl_types.all;
entity keyboard1_tb is
end keyboard1_tb;
