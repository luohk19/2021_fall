library verilog;
use verilog.vl_types.all;
entity MyClock_vlg_check_tst is
    port(
        num0            : in     vl_logic;
        num1            : in     vl_logic;
        num2            : in     vl_logic;
        num3            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end MyClock_vlg_check_tst;
