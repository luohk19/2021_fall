library verilog;
use verilog.vl_types.all;
entity MyClock_vlg_vec_tst is
end MyClock_vlg_vec_tst;
